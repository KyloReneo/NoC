-- THE TOP LEVEL MODULE OF THE ROUTER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY ROUTER IS
	GENERIC(
		NODE_ADDRESS : NETWORK_ADDR
	);
	PORT(
		-- GLOBAL CLOCK AND RESET SIGNALS
        	CLK               : IN STD_LOGIC;
        	RST               : IN STD_LOGIC;
		-- HANDLING INPUT BUFFERS
		-- INPUT PORTS FOR ADJACENT ROUTERS
        	NORTH_DATA_IN     : IN FLIT;
        	EAST_DATA_IN      : IN FLIT;
        	SOUTH_DATA_IN     : IN FLIT;
        	WEST_DATA_IN      : IN FLIT;
		-- PORTS FOR CHECKING CREDIT OUT OF ADJACENT BUFFERS
        	NORTH_CREDIT_IN   : IN STD_LOGIC;
        	EAST_CREDIT_IN    : IN STD_LOGIC;
        	SOUTH_CREDIT_IN   : IN STD_LOGIC;
        	WEST_CREDIT_IN    : IN STD_LOGIC;
		-- WRITE REQUEST SIGNALS COMES FROM ADJACENT ROUTERS
        	NORTH_WR_REQ_IN   : IN STD_LOGIC;
        	EAST_WR_REQ_IN    : IN STD_LOGIC;
        	SOUTH_WR_REQ_IN   : IN STD_LOGIC;
        	WEST_WR_REQ_IN    : IN STD_LOGIC;
		-- OUTPUT PORTS TO ADJACENT ROUTERS 
		LOCAL_DATA_OUT    : OUT FLIT;
        	NORTH_DATA_OUT    : OUT FLIT;
        	EAST_DATA_OUT     : OUT FLIT;
        	SOUTH_DATA_OUT    : OUT FLIT;
        	WEST_DATA_OUT     : OUT FLIT;
		-- ROUTER'S OUTPUT SIGNALS
		LOCAL_CREDIT_OUT  : OUT STD_LOGIC;
        	NORTH_CREDIT_OUT  : OUT STD_LOGIC;
        	EAST_CREDIT_OUT   : OUT STD_LOGIC;
        	SOUTH_CREDIT_OUT  : OUT STD_LOGIC;
        	WEST_CREDIT_OUT   : OUT STD_LOGIC;
		-- WRITE REQUEST SIGNALS TO ADJACENT ROUTERS
        	NORTH_WR_REQ_OUT  : OUT STD_LOGIC;
        	EAST_WR_REQ_OUT   : OUT STD_LOGIC;
        	SOUTH_WR_REQ_OUT  : OUT STD_LOGIC;
        	WEST_WR_REQ_OUT   : OUT STD_LOGIC;
		-- IP CORE RELATED INPUT AND OUTPUTS
        	-- NI SIDE FORM THE INJECTOR CHANNEL
		FLIT_DEST_ADDR_TO_NI : IN    NETWORK_ADDR;
		HEAD_OR_TAIL         : IN    STD_LOGIC;
        	VALID_TO_NI          : IN    STD_LOGIC;
		READY_FROM_NI        : OUT   STD_LOGIC;
        	-- NI SIDE FORM THE EXTRACTOR CHANNEL  
		READY_TO_NI          : IN    STD_LOGIC;                                    -- IP CORE IS READY TO RECEIVE DATA FROM NI
        	PAYLOAD_FORM_NI      : OUT   STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0); -- FOR THIS PROJECT WE ASSUME THAT THE PAYLOAD IS SOURCE ADDRESS OF THE FLIT THAT RECEIVED AT THE NI EXTRACTOR CHANNEL OK?!
        	VALID_FROM_NI        : OUT   STD_LOGIC                                     -- DATA IN NI IS READY
        	
	);

END ENTITY ROUTER;

ARCHITECTURE STRUCT OF ROUTER IS

-- COMPONENT DECLRATIONS
-- INPUT BUFFER COMPONENT
COMPONENT INPUT_BUFFER
	PORT(
		CLK 	           : IN  STD_LOGIC;
		RST	           : IN  STD_LOGIC;
		WRITE_REQUEST      : IN  STD_LOGIC;
		GRANT  	           : IN  STD_LOGIC;
		CREDIT_IN          : IN  STD_LOGIC; 					
		DATA               : IN  FLIT;
		REQUEST_TO_ARBITER : OUT NETWORK_ADDR;
		CREDIT_OUT         : OUT STD_LOGIC; 					
		EMPTY              : OUT STD_LOGIC;
		OUTPUT             : OUT FLIT
		);
END COMPONENT;
-- EXTRACTOR BUFFER COMPONENT
COMPONENT EXTRACTOR_BUFFER
	PORT(
		CLK 	           : IN  STD_LOGIC;
		RST	           : IN  STD_LOGIC;
		WRITE_REQUEST      : IN  STD_LOGIC;
		GRANT  	           : IN  STD_LOGIC;
		DATA               : IN  FLIT;
		CREDIT_OUT         : OUT STD_LOGIC; 					
		EMPTY              : OUT STD_LOGIC;
		OUTPUT             : OUT FLIT
		);
END COMPONENT;
-- CROSSBAR SWITCH COMPONENT
COMPONENT CROSSBAR_SWITCH
    PORT (
        DATA_LOCAL_IN  : IN  FLIT;  
        DATA_NORTH_IN  : IN  FLIT;
        DATA_EAST_IN   : IN  FLIT;
        DATA_SOUTH_IN  : IN  FLIT;
        DATA_WEST_IN   : IN  FLIT; 
        SEL_LOCAL      : IN  DIRECTION; 
        SEL_NORTH      : IN  DIRECTION;
        SEL_EAST       : IN  DIRECTION;
        SEL_SOUTH      : IN  DIRECTION;
        SEL_WEST       : IN  DIRECTION;
        DATA_LOCAL_OUT : OUT FLIT;
        DATA_NORTH_OUT : OUT FLIT;
        DATA_EAST_OUT  : OUT FLIT;
        DATA_SOUTH_OUT : OUT FLIT;
        DATA_WEST_OUT  : OUT FLIT  
    );
END COMPONENT;
-- ARBITER COMPONENT
COMPONENT ARBITER
    PORT (
        CLK                 : IN STD_LOGIC;
        RST                 : IN STD_LOGIC;
        -- EMPTY FLAGS FROM INPUT BUFFERS (ACTIVE HIGH '1' MEANS EMPTY, '0' MEANS HAS DATA)
        EMPTY_IN_LOCAL      : IN STD_LOGIC;
        EMPTY_IN_NORTH      : IN STD_LOGIC;
        EMPTY_IN_EAST       : IN STD_LOGIC;
        EMPTY_IN_SOUTH      : IN STD_LOGIC;
        EMPTY_IN_WEST       : IN STD_LOGIC;
        -- DESTINATION ADDRESSES FROM INPUT BUFFERS (THE HEAD FLIT OF EACH FIFO)
        DEST_ADDR_IN_LOCAL  : IN NETWORK_ADDR;
        DEST_ADDR_IN_NORTH  : IN NETWORK_ADDR;
        DEST_ADDR_IN_EAST   : IN NETWORK_ADDR;
        DEST_ADDR_IN_SOUTH  : IN NETWORK_ADDR;
        DEST_ADDR_IN_WEST   : IN NETWORK_ADDR;
        -- OUTPUTS TO ROUTING UNITS (THE DESTINATION ADDRESSES TO BE ROUTED)
        DEST_ADDR_OUT_LOCAL : OUT NETWORK_ADDR;
        DEST_ADDR_OUT_NORTH : OUT NETWORK_ADDR;
        DEST_ADDR_OUT_EAST  : OUT NETWORK_ADDR;
        DEST_ADDR_OUT_SOUTH : OUT NETWORK_ADDR;
        DEST_ADDR_OUT_WEST  : OUT NETWORK_ADDR;
        -- INPUTS FROM ROUTING UNITS (THE CALCULATED OUTPUT DIRECTION FOR EACH INPUT)
        ROUTE_DIR_IN_LOCAL  : IN DIRECTION;
        ROUTE_DIR_IN_NORTH  : IN DIRECTION;
        ROUTE_DIR_IN_EAST   : IN DIRECTION;
        ROUTE_DIR_IN_SOUTH  : IN DIRECTION;
        ROUTE_DIR_IN_WEST   : IN DIRECTION;
        -- GRANTS TO INPUT BUFFERS (READ ENABLE SIGNALS)
        GRANT_OUT_LOCAL     : OUT STD_LOGIC;
        GRANT_OUT_NORTH     : OUT STD_LOGIC;
        GRANT_OUT_EAST      : OUT STD_LOGIC;
        GRANT_OUT_SOUTH     : OUT STD_LOGIC;
        GRANT_OUT_WEST      : OUT STD_LOGIC;
        -- CREDIT-BASED FLOW CONTROL FROM DOWNSTREAM ROUTERS
        -- '0' MEANS THE ADJASENT INPUT BUFFER IS NOT FULL (CREDIT AVAILABLE)
        CREDIT_IN_LOCAL     : IN STD_LOGIC;
        CREDIT_IN_NORTH     : IN STD_LOGIC;
        CREDIT_IN_EAST      : IN STD_LOGIC;
        CREDIT_IN_SOUTH     : IN STD_LOGIC;
        CREDIT_IN_WEST      : IN STD_LOGIC;
        -- WRITE REQUEST TO TARGET BUFFERS IN THE NEXT ROUTER
        W_REQ_OUT_LOCAL     : OUT STD_LOGIC;
        W_REQ_OUT_NORTH     : OUT STD_LOGIC;
        W_REQ_OUT_EAST      : OUT STD_LOGIC;
        W_REQ_OUT_SOUTH     : OUT STD_LOGIC;
        W_REQ_OUT_WEST      : OUT STD_LOGIC;
        -- SELECT SIGNALS FOR THE 5 OUTPUT CROSSBARS (ONE PER OUTPUT PORT)
        SEL_LOCAL           : OUT DIRECTION; 
        SEL_NORTH           : OUT DIRECTION;
        SEL_EAST            : OUT DIRECTION;
        SEL_SOUTH           : OUT DIRECTION;
        SEL_WEST            : OUT DIRECTION;
	-- CREDIT OUT TO THE GRANTED INPUT BUFFER
	CREDIT_OUT          : OUT STD_LOGIC
    );
END COMPONENT;
-- ROUTING UNIT COMPONENT
COMPONENT ROUTING_UNIT
     GENERIC(
	NODE_ADDRESS : NETWORK_ADDR
    );
    PORT (
        DEST_ADDRESS : IN  NETWORK_ADDR; -- THE DESTINATION PART OF EACH HEADER FLIT COMES FROM THE FIFO BUFFER
        ROUTE_DIR    : OUT DIRECTION     -- THE REQUESTED OUTPUT DIRECTION
    );
END COMPONENT;
--NETWORK INTERFACE COMPONENT
COMPONENT NETWORK_INTERFACE
    GENERIC (
        NODE_ADDR  : NETWORK_ADDR
    );
    PORT (
        CLK                     : IN STD_LOGIC;
        RST                     : IN STD_LOGIC;

        -- IP CORE SIDE
	-- TO INJECTOR CHANNEL
        FLIT_DEST_ADDR_FORM_IP  : IN  NETWORK_ADDR;
	HEAD_OR_TAIL            : IN  STD_LOGIC;
        VALID_IN_FROM_IP        : IN  STD_LOGIC;
        READY_OUT_TO_IP         : OUT STD_LOGIC;
	-- FROM EXTRACTOR CHANNEL
	READY_FROM_IP           : IN  STD_LOGIC;
	VALID_TO_IP             : OUT STD_LOGIC;
        PAYLOAD_TO_IP           : OUT STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        -- ROUTER SIDE 
        -- TO ROUTER'S LOCAL INPUT BUFFER (BUFFERED OUTPUT)
        LOCAL_IB_FULL   : IN  STD_LOGIC;  -- LOCAL INPUT BUFFER'S FULL FLAG
	LOCAL_IB_WR     : OUT STD_LOGIC;  -- WRITE ENABLE SIGNAL TO LOCAL INPUT BUFFER
        LOCAL_IB_DATA   : OUT FLIT;       -- DATA TO LOCAL INPUT BUFFER
        -- FROM ROUTER'S CROSSBAR TO EXTRACTOR CHANNEL (UNBUFFERED OUTPUT OF ROUTER)
        ROUTER_TO_NI    : IN  FLIT;       -- DIRECTLY COMES FROM CROSSBAR OUTPUT
	-- CONTROLLING SIGNALS TO AND FROM ARBITTER FOR THE EXTRACTOR CHANNEL
	EXT_W_REQ_IN   : IN  STD_LOGIC;
	EXT_CREDIT_OUT : OUT STD_LOGIC
        -- noc_ext_valid   : IN  STD_LOGIC;  -- Crossbar has valid data for us
        -- noc_ext_ready   : OUT STD_LOGIC   -- NI IS READY TO ACCEPT THE DATA 
    );
END COMPONENT;

-- INTERNAL CONNECTIONS AND SIGNALS
-- INPUT BUFFERS INTERCONNECTIONS (OUTPUTS)
SIGNAL LOCAL_IB_DATA,       NORTH_IB_DATA,       EAST_IB_DATA,       SOUTH_IB_DATA,       WEST_IB_DATA       : FLIT;
SIGNAL LOCAL_IB_EMPTY,      NORTH_IB_EMPTY,      EAST_IB_EMPTY,      SOUTH_IB_EMPTY,      WEST_IB_EMPTY      : STD_LOGIC;
SIGNAL LOCAL_IB_CREDIT_OUT, NORTH_IB_CREDIT_OUT, EAST_IB_CREDIT_OUT, SOUTH_IB_CREDIT_OUT, WEST_IB_CREDIT_OUT : STD_LOGIC;


-- CREDIT SIGNAL BETWEEN ARBITER AND EXTRACTOR CHANNEL
SIGNAL LOCAL_IB_CREDIT_IN : STD_LOGIC;

-- ARBITER INTERCONNECTIONS (OUTPUTS)    
SIGNAL ARB_GRANT_LOCAL,  ARB_GRANT_NORTH,  ARB_GRANT_EAST,  ARB_GRANT_SOUTH,  ARB_GRANT_WEST  : STD_LOGIC;
SIGNAL ARB_WR_REQ_LOCAL, ARB_WR_REQ_NORTH, ARB_WR_REQ_EAST, ARB_WR_REQ_SOUTH, ARB_WR_REQ_WEST : STD_LOGIC;    
SIGNAL ARB_SEL_LOCAL,    ARB_SEL_NORTH,    ARB_SEL_EAST,    ARB_SEL_SOUTH,    ARB_SEL_WEST    : DIRECTION;
SIGNAL ARB_TO_IB_CREDIT : STD_LOGIC;

-- CROSSBAR INTERCONNECTIONS (OUTPUTS)    
SIGNAL XBAR_OUT_LOCAL, XBAR_OUT_NORTH, XBAR_OUT_EAST, XBAR_OUT_SOUTH, XBAR_OUT_WEST : FLIT;

-- ROUTING UNITS INTERCONNECTIONS (OUTPUTS)    
SIGNAL ROUTING_DEST_LOCAL, ROUTING_DEST_NORTH, ROUTING_DEST_EAST, ROUTING_DEST_SOUTH, ROUTING_DEST_WEST : NETWORK_ADDR;
SIGNAL RU_DEST_LOCAL, RU_DEST_NORTH, RU_DEST_EAST, RU_DEST_SOUTH, RU_DEST_WEST                          : NETWORK_ADDR;
SIGNAL ROUTING_DIR_LOCAL,  ROUTING_DIR_NORTH,  ROUTING_DIR_EAST,  ROUTING_DIR_SOUTH,  ROUTING_DIR_WEST  : DIRECTION;
    
-- NI AND IP CORE SIGNALS
SIGNAL NI_TO_LOCAL_WR, NI_TO_LOCAL_FULL : STD_LOGIC;
SIGNAL NI_TO_LOCAL_DATA                 : FLIT;

-- IP CORE RELATED SIGNALS
SIGNAL RFNI, VFNI : STD_LOGIC;
SIGNAL PFNI : NETWORK_ADDR;

BEGIN

-- COMPONRNT INSTANTIATION
-- INPUT BUFFERS FOR EACH DIRECTION
    LOCAL_INPUT_BUFFER : INPUT_BUFFER
        PORT MAP(
            CLK                 => CLK,
            RST                 => RST,
            WRITE_REQUEST       => NI_TO_LOCAL_WR,
	    GRANT  	        => ARB_GRANT_LOCAL,
	    CREDIT_IN           => ARB_TO_IB_CREDIT,					
	    DATA                => NI_TO_LOCAL_DATA,
	    REQUEST_TO_ARBITER  => ROUTING_DEST_LOCAL,
	    CREDIT_OUT          => LOCAL_IB_CREDIT_OUT,					
	    EMPTY               => LOCAL_IB_EMPTY,
	    OUTPUT		=> LOCAL_IB_DATA
        );
    NORTH_INPUT_BUFFER : INPUT_BUFFER
        PORT MAP(
            CLK                 => CLK,
            RST                 => RST,
            WRITE_REQUEST       => NORTH_WR_REQ_IN,
	    GRANT  	        => ARB_GRANT_NORTH,
	    CREDIT_IN           => ARB_TO_IB_CREDIT,					
	    DATA                => NORTH_DATA_IN,
	    REQUEST_TO_ARBITER  => ROUTING_DEST_NORTH,
	    CREDIT_OUT          => NORTH_IB_CREDIT_OUT,					
	    EMPTY               => NORTH_IB_EMPTY,
	    OUTPUT		=> NORTH_IB_DATA
        );
    EAST_INPUT_BUFFER : INPUT_BUFFER
        PORT MAP(
            CLK                 => CLK,
            RST                 => RST,
            WRITE_REQUEST       => EAST_WR_REQ_IN,
	    GRANT  	        => ARB_GRANT_EAST,
	    CREDIT_IN           => ARB_TO_IB_CREDIT,					
	    DATA                => EAST_DATA_IN,
	    REQUEST_TO_ARBITER  => ROUTING_DEST_EAST,
	    CREDIT_OUT          => EAST_IB_CREDIT_OUT,					
	    EMPTY               => EAST_IB_EMPTY,
	    OUTPUT		=> EAST_IB_DATA
        );
    SOUTH_INPUT_BUFFER : INPUT_BUFFER
        PORT MAP(
            CLK                 => CLK,
            RST                 => RST,
            WRITE_REQUEST       => SOUTH_WR_REQ_IN,
	    GRANT  	        => ARB_GRANT_SOUTH,
	    CREDIT_IN           => ARB_TO_IB_CREDIT,					
	    DATA                => SOUTH_DATA_IN,
	    REQUEST_TO_ARBITER  => ROUTING_DEST_SOUTH,
	    CREDIT_OUT          => SOUTH_IB_CREDIT_OUT,					
	    EMPTY               => SOUTH_IB_EMPTY,
	    OUTPUT		=> SOUTH_IB_DATA
        );
    WEST_INPUT_BUFFER : INPUT_BUFFER
        PORT MAP(
            CLK                 => CLK,
            RST                 => RST,
            WRITE_REQUEST       => WEST_WR_REQ_IN,
	    GRANT  	        => ARB_GRANT_WEST,
	    CREDIT_IN           => ARB_TO_IB_CREDIT,					
	    DATA                => WEST_DATA_IN,
	    REQUEST_TO_ARBITER  => ROUTING_DEST_WEST,
	    CREDIT_OUT          => WEST_IB_CREDIT_OUT,					
	    EMPTY               => WEST_IB_EMPTY,
	    OUTPUT		=> WEST_IB_DATA
        );
-- ROUTING UNITS FOR EACH INPUT BUFFER
    LOCAL_ROUTING_UNIT : ROUTING_UNIT
	GENERIC MAP(
	NODE_ADDRESS            => NODE_ADDRESS
        )
        PORT MAP(
            DEST_ADDRESS        => RU_DEST_LOCAL,
            ROUTE_DIR           => ROUTING_DIR_LOCAL
        );
    NORTH_ROUTING_UNIT : ROUTING_UNIT
	GENERIC MAP(
	NODE_ADDRESS            => NODE_ADDRESS
        )
        PORT MAP(
            DEST_ADDRESS        => RU_DEST_NORTH,
            ROUTE_DIR           => ROUTING_DIR_NORTH
        );
    EAST_ROUTING_UNIT  : ROUTING_UNIT
	GENERIC MAP(
	NODE_ADDRESS            => NODE_ADDRESS
        )
        PORT MAP(
            DEST_ADDRESS        => RU_DEST_EAST,
            ROUTE_DIR           => ROUTING_DIR_EAST
        );
    SOUTH_ROUTING_UNIT : ROUTING_UNIT
	GENERIC MAP(
	NODE_ADDRESS            => NODE_ADDRESS
        )
        PORT MAP(
            DEST_ADDRESS        => RU_DEST_SOUTH,
            ROUTE_DIR           => ROUTING_DIR_SOUTH
        );
    WEST_ROUTING_UNIT  : ROUTING_UNIT
	GENERIC MAP(
	NODE_ADDRESS            => NODE_ADDRESS
        )
        PORT MAP(
            DEST_ADDRESS        => RU_DEST_WEST,
            ROUTE_DIR           => ROUTING_DIR_WEST
        ); 
-- ARBITER
   ROUTER_ARBITER : ARBITER
	PORT MAP(
	    CLK  		=> CLK,
            RST 		=> RST,
            EMPTY_IN_LOCAL 	=> LOCAL_IB_EMPTY,
            EMPTY_IN_NORTH 	=> NORTH_IB_EMPTY,
            EMPTY_IN_EAST  	=> EAST_IB_EMPTY,
            EMPTY_IN_SOUTH 	=> SOUTH_IB_EMPTY,
            EMPTY_IN_WEST  	=> WEST_IB_EMPTY,
            DEST_ADDR_IN_LOCAL  => ROUTING_DEST_LOCAL,
            DEST_ADDR_IN_NORTH  => ROUTING_DEST_NORTH,
            DEST_ADDR_IN_EAST   => ROUTING_DEST_EAST,
            DEST_ADDR_IN_SOUTH  => ROUTING_DEST_SOUTH,
            DEST_ADDR_IN_WEST   => ROUTING_DEST_WEST,
            DEST_ADDR_OUT_LOCAL => RU_DEST_LOCAL,
            DEST_ADDR_OUT_NORTH => RU_DEST_NORTH,
            DEST_ADDR_OUT_EAST  => RU_DEST_EAST,
            DEST_ADDR_OUT_SOUTH => RU_DEST_SOUTH,
            DEST_ADDR_OUT_WEST  => RU_DEST_WEST,
            ROUTE_DIR_IN_LOCAL  => ROUTING_DIR_LOCAL,
            ROUTE_DIR_IN_NORTH  => ROUTING_DIR_NORTH,
            ROUTE_DIR_IN_EAST   => ROUTING_DIR_EAST,
            ROUTE_DIR_IN_SOUTH  => ROUTING_DIR_SOUTH,
            ROUTE_DIR_IN_WEST   => ROUTING_DIR_WEST,
            GRANT_OUT_LOCAL     => ARB_GRANT_LOCAL,
            GRANT_OUT_NORTH     => ARB_GRANT_NORTH,
            GRANT_OUT_EAST      => ARB_GRANT_EAST,
            GRANT_OUT_SOUTH     => ARB_GRANT_SOUTH,
            GRANT_OUT_WEST      => ARB_GRANT_WEST,
            CREDIT_IN_LOCAL     => LOCAL_IB_CREDIT_IN, -- CREDIT_OUT THAT COMES FROM EXTRACTOR CHANNEL
            CREDIT_IN_NORTH     => NORTH_CREDIT_IN,
            CREDIT_IN_EAST      => EAST_CREDIT_IN,
            CREDIT_IN_SOUTH     => SOUTH_CREDIT_IN,
            CREDIT_IN_WEST      => WEST_CREDIT_IN,
            W_REQ_OUT_LOCAL     => ARB_WR_REQ_LOCAL,
            W_REQ_OUT_NORTH     => ARB_WR_REQ_NORTH,
            W_REQ_OUT_EAST      => ARB_WR_REQ_EAST,
            W_REQ_OUT_SOUTH     => ARB_WR_REQ_SOUTH,
            W_REQ_OUT_WEST      => ARB_WR_REQ_WEST,
            SEL_LOCAL 		=> ARB_SEL_LOCAL,
            SEL_NORTH 		=> ARB_SEL_NORTH,
            SEL_EAST  		=> ARB_SEL_EAST,
            SEL_SOUTH 		=> ARB_SEL_SOUTH,
            SEL_WEST  		=> ARB_SEL_WEST,
	    CREDIT_OUT          => ARB_TO_IB_CREDIT
	);
-- CROSSBAR SWITCH
   CROSSBAR : CROSSBAR_SWITCH
	PORT MAP(
	    DATA_LOCAL_IN  	=> LOCAL_IB_DATA,
            DATA_NORTH_IN 	=> NORTH_IB_DATA,
            DATA_EAST_IN   	=> EAST_IB_DATA,
            DATA_SOUTH_IN  	=> SOUTH_IB_DATA,
            DATA_WEST_IN   	=> WEST_IB_DATA, 
            SEL_LOCAL      	=> ARB_SEL_LOCAL,
            SEL_NORTH      	=> ARB_SEL_NORTH,
            SEL_EAST       	=> ARB_SEL_EAST,
            SEL_SOUTH      	=> ARB_SEL_SOUTH,
            SEL_WEST       	=> ARB_SEL_WEST,
            DATA_LOCAL_OUT 	=> XBAR_OUT_LOCAL,
            DATA_NORTH_OUT 	=> XBAR_OUT_NORTH,
            DATA_EAST_OUT  	=> XBAR_OUT_EAST,
            DATA_SOUTH_OUT 	=> XBAR_OUT_SOUTH,
            DATA_WEST_OUT  	=> XBAR_OUT_WEST
	);
-- NETWORK INTERFACE
   NI      : NETWORK_INTERFACE
	GENERIC MAP(
             NODE_ADDR  => NODE_ADDRESS
    	)
	PORT MAP(
	    CLK                     => CLK,
            RST                     => RST,
            FLIT_DEST_ADDR_FORM_IP  => FLIT_DEST_ADDR_TO_NI,
	    HEAD_OR_TAIL            => HEAD_OR_TAIL,
            VALID_IN_FROM_IP        => VALID_TO_NI,
            READY_OUT_TO_IP         => RFNI,
	    READY_FROM_IP           => READY_TO_NI,
	    VALID_TO_IP             => VFNI,
            PAYLOAD_TO_IP           => PFNI,
            LOCAL_IB_FULL   	    => LOCAL_IB_CREDIT_OUT,
	    LOCAL_IB_WR     	    => NI_TO_LOCAL_WR,
            LOCAL_IB_DATA   	    => NI_TO_LOCAL_DATA,
            ROUTER_TO_NI    	    => XBAR_OUT_LOCAL,
	    EXT_W_REQ_IN    	    => ARB_WR_REQ_LOCAL,
	    EXT_CREDIT_OUT          => LOCAL_IB_CREDIT_IN   -- EXTRACTOR BUFFER FULL FLAG
	);

 -- OUTPUT PORTS CONNECTIONS
    LOCAL_DATA_OUT <= XBAR_OUT_LOCAL;
    NORTH_DATA_OUT <= XBAR_OUT_NORTH;
    EAST_DATA_OUT  <= XBAR_OUT_EAST;
    SOUTH_DATA_OUT <= XBAR_OUT_SOUTH;
    WEST_DATA_OUT  <= XBAR_OUT_WEST;

    -- CREDIT OUT SIGNALS
    LOCAL_CREDIT_OUT <= LOCAL_IB_CREDIT_OUT;
    NORTH_CREDIT_OUT <= NORTH_IB_CREDIT_OUT;
    EAST_CREDIT_OUT  <= EAST_IB_CREDIT_OUT;
    SOUTH_CREDIT_OUT <= SOUTH_IB_CREDIT_OUT;
    WEST_CREDIT_OUT  <= WEST_IB_CREDIT_OUT;

    -- WRITE REQUEST OUTPUTS
    NORTH_WR_REQ_OUT <= ARB_WR_REQ_NORTH;
    EAST_WR_REQ_OUT  <= ARB_WR_REQ_EAST;
    SOUTH_WR_REQ_OUT <= ARB_WR_REQ_SOUTH;
    WEST_WR_REQ_OUT  <= ARB_WR_REQ_WEST;

    -- IP CORE 
    READY_FROM_NI    <= RFNI;
    PAYLOAD_FORM_NI  <= PFNI;
    VALID_FROM_NI    <= VFNI;

END ARCHITECTURE STRUCT;
