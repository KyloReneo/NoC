-- SINGLE ROUTING UNIT (WE HAVE TO DEDICATE A ROUTING UNIT TO EACH INPUT BUFFER FOR THE BETTER EXPERIENCE, SO WE NEED 5 OF THIS IN THE TOP LEVEL MODULE)
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY ROUTING_UNIT IS
    GENERIC(
	NODE_ADDRESS : NETWORK_ADDR
    );
    PORT (
        DEST_ADDRESS : IN  NETWORK_ADDR; -- THE DESTINATION PART OF EACH HEADER FLIT COMES FROM THE FIFO BUFFER
        ROUTE_DIR    : OUT DIRECTION     -- THE REQUESTED OUTPUT DIRECTION
    );
END ENTITY;

ARCHITECTURE BEHAV OF ROUTING_UNIT IS
    SIGNAL DESTINATION_X, DESTINATION_Y : INTEGER;
    SIGNAL CURRENT_X,     CURRENT_Y     : INTEGER;
    BEGIN
    -- DESTINATION COORDINATES
    DESTINATION_X <= ADDRESS_X(DEST_ADDRESS);
    DESTINATION_Y <= ADDRESS_Y(DEST_ADDRESS);
    CURRENT_X     <= ADDRESS_X(NODE_ADDRESS);
    CURRENT_Y     <= ADDRESS_Y(NODE_ADDRESS);

    -- XY Routing Algorithm Process
    PROCESS(DESTINATION_X, DESTINATION_Y, CURRENT_X, CURRENT_Y)
    BEGIN
        ROUTE_DIR <= DISCONNECTED;

        -- ROUTE IN X DIRECTION FIRST, THEN ROUTE IN Y DIRECTION AND IF BOTH X & Y ARE EQUAL CURRENT NODE IS THE DESTINATION
        IF    CURRENT_X < DESTINATION_X THEN
            ROUTE_DIR <= EAST;
        ELSIF CURRENT_X > DESTINATION_X THEN
            ROUTE_DIR <= WEST;
        ELSIF CURRENT_Y < DESTINATION_Y THEN
            ROUTE_DIR <= SOUTH;
        ELSIF CURRENT_Y > DESTINATION_Y THEN
            ROUTE_DIR <= NORTH;
        ELSE
            ROUTE_DIR <= LOCAL;
        END IF;
    END PROCESS;
END ARCHITECTURE BEHAV;
