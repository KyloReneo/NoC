-- MULTIPLEXR USED IN CROSSBAR SWITCH
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY CROSSBAR_MUX_EAST IS
    PORT (
        LOCAL_IN : IN  FLIT;
        NORTH_IN : IN  FLIT;
        SOUTH_IN : IN  FLIT;
        WEST_IN  : IN  FLIT;
        SEL      : IN  DIRECTION;
        DATA_OUT : OUT FLIT
    );
END ENTITY;

ARCHITECTURE BEHAV OF CROSSBAR_MUX_EAST IS
BEGIN
    WITH SEL SELECT DATA_OUT <=
        LOCAL_IN WHEN LOCAL,
        NORTH_IN WHEN NORTH,
        SOUTH_IN WHEN SOUTH,
        WEST_IN  WHEN WEST,
        (OTHERS => '0') WHEN OTHERS;
END ARCHITECTURE;
