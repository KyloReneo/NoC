-- PACKAGE FOR COMMON TYPES AND CONSTANTS
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE ROUTER_PKG IS

-- NETWORK ADDRESS PARAMS
CONSTANT DATA_WIDTH        : INTEGER := 12;
CONSTANT FLIT_TYPE_WIDTH   : INTEGER := 2;
CONSTANT ADDRESS_WIDTH     : INTEGER := 5; -- NETWORK ADDRESS WIDTH

-- SUBTYPES
SUBTYPE NETWORK_ADDR IS STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
SUBTYPE FLIT         IS STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);

-- NODE ADDRESS
CONSTANT NODE5_ADDRESS : NETWORK_ADDR := "00101"; -- THIS IS NODE 5
CONSTANT NODE6_ADDRESS : NETWORK_ADDR := "00110"; -- THIS IS NODE 6

-- TOPOLOGY INFO
CONSTANT ROWS    : INTEGER := 4;
CONSTANT COLUMNS : INTEGER := 4;


-- FIFO BUFFER RELATED CONSTANTS
CONSTANT BUFFER_DEPTH      : INTEGER := 8;
CONSTANT BUFFER_PTR_WIDTH  : INTEGER := 3;

-- ARBITER

-- XBAR
CONSTANT XBAR_KEY_SIZE : INTEGER := 2;
CONSTANT MUX_ADDR_BIT  : INTEGER := 3; -- HOW MANY BITS NEEDED TO ADDRESSING ALL MULTIPLEXERS IN THE CROSSBAR

-- PHYSICAL DIRECTIONS OF EACH ROUTER
TYPE DIRECTION IS (LOCAL, NORTH, EAST, SOUTH, WEST, DISCONNECTED);

-- FUNCTIONS
FUNCTION ADDRESS_X(FLIT_DESTINATION : NETWORK_ADDR) RETURN INTEGER;
FUNCTION ADDRESS_Y(FLIT_DESTINATION : NETWORK_ADDR) RETURN INTEGER;

END PACKAGE;

PACKAGE BODY ROUTER_PKG IS
-- A FUNCTION TO RETURN THE X OF THE DESTINATION OF THE FLITS COMMING FROM THE ARBITER
FUNCTION ADDRESS_X(FLIT_DESTINATION : NETWORK_ADDR) RETURN INTEGER IS
    BEGIN
        RETURN TO_INTEGER(UNSIGNED(FLIT_DESTINATION(ADDRESS_WIDTH - 1 DOWNTO 0))) MOD COLUMNS;
END FUNCTION;
-- A FUNCTION TO RETURN THE X OF THE DESTINATION OF THE FLITS COMMING FROM THE ARBITER
FUNCTION ADDRESS_Y(FLIT_DESTINATION : NETWORK_ADDR) RETURN INTEGER IS
    BEGIN
        RETURN TO_INTEGER(UNSIGNED(FLIT_DESTINATION(ADDRESS_WIDTH - 1 DOWNTO 0))) / ROWS;
END FUNCTION;

END PACKAGE BODY;
