-- MULTIPLEXR USED IN CROSSBAR SWITCH
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY CROSSBAR_MUX_WEST IS
    PORT (
        LOCAL_IN : IN  FLIT;
        NORTH_IN : IN  FLIT;
        EAST_IN  : IN  FLIT;
        SOUTH_IN : IN  FLIT;
        SEL      : IN  DIRECTION;
        DATA_OUT : OUT FLIT
    );
END ENTITY;

ARCHITECTURE BEHAV OF CROSSBAR_MUX_WEST IS
BEGIN
    WITH SEL SELECT DATA_OUT <=
        LOCAL_IN WHEN LOCAL,
        NORTH_IN WHEN NORTH,
        EAST_IN  WHEN EAST,
        SOUTH_IN WHEN SOUTH,
        (OTHERS => '0') WHEN OTHERS;
END ARCHITECTURE;
