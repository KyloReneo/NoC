-- A CONFIGURABLE EXTRACTOR BUFFER OF THE NETWORK INTERFACE OF EACH ROUTER THAT GETS DATA FROM ADJASENT ROUTERS AND SENDS IT TO IP CORE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY EXTRACTOR_BUFFER IS
	PORT(
		CLK 	           : IN  STD_LOGIC;
		RST	           : IN  STD_LOGIC;
		WRITE_REQUEST      : IN  STD_LOGIC;
		GRANT  	           : IN  STD_LOGIC;
		IP_REQ		   : IN  STD_LOGIC;
		DATA               : IN  FLIT;
		CREDIT_OUT         : OUT STD_LOGIC; 					
		EMPTY              : OUT STD_LOGIC;
		OUTPUT             : OUT FLIT
		);
END EXTRACTOR_BUFFER;

ARCHITECTURE BEHAV OF EXTRACTOR_BUFFER IS

-- COMPONENTS DECLARATIONS
-- FIFO CONTROLLER
COMPONENT FIFO_CONTROLLER 
	PORT(
		FC_CLK   : IN  STD_LOGIC;
		FC_RST   : IN  STD_LOGIC;
		FC_WR    : IN  STD_LOGIC;
		FC_RD    : IN  STD_LOGIC;
		FC_FULL  : OUT STD_LOGIC;
		FC_EMPTY : OUT STD_LOGIC;
		WR_EN    : OUT STD_LOGIC;
		WR_ADDR  : OUT STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0);
		RE_ADDR  : OUT STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0)
		);
END COMPONENT;

-- REGISTER FILE
COMPONENT REGISTER_FILE 
    PORT (
        RF_CLK             : IN  STD_LOGIC;
	RF_RST             : IN  STD_LOGIC;
        WR_EN              : IN  STD_LOGIC;
	GRANT              : IN  STD_LOGIC;
	CREDIT_IN          : IN  STD_LOGIC;
	EMPTY              : IN  STD_LOGIC;
        WR_ADDR            : IN  STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0);
        RE_ADDR            : IN  STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0);
        DATA_IN            : IN  STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
	REQUEST_TO_ARBITER : OUT STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        DATA_OUT           : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
    	);
END COMPONENT;

-- INTERNAL CONNECTIONS
SIGNAL REG_WRITE_EN  : STD_LOGIC;
SIGNAL W_ADDR        : STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0) := (OTHERS => '1');
SIGNAL R_ADDR        : STD_LOGIC_VECTOR(BUFFER_PTR_WIDTH - 1 DOWNTO 0) := (OTHERS => '1');

BEGIN



-- COMPONENTS INSTANTIATIONS
-- FIFO CONTROLLER
CONTROLLER_INST : FIFO_CONTROLLER 
	PORT MAP(
		FC_CLK   => CLK,
		FC_RST   => RST,
		FC_WR    => WRITE_REQUEST,
		FC_RD    => GRANT,
		FC_FULL  => CREDIT_OUT,
		FC_EMPTY => EMPTY,
		WR_EN    => REG_WRITE_EN,
		WR_ADDR  => W_ADDR,
		RE_ADDR  => R_ADDR
		);

-- REGISTER FILE
RF_INST : REGISTER_FILE 
	PORT MAP(
        	RF_CLK             => CLK,
		RF_RST             => RST,
        	WR_EN              => REG_WRITE_EN,
		GRANT              => GRANT,
		CREDIT_IN          => IP_REQ,
		EMPTY              => EMPTY,
        	WR_ADDR            => W_ADDR,
        	RE_ADDR            => R_ADDR,
        	DATA_IN            => DATA,
		REQUEST_TO_ARBITER => OPEN,
        	DATA_OUT           => OUTPUT
    		);
END BEHAV;
