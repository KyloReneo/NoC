-- ROUTERS 5 AND 6 OF THE 4*4 MESH CONNECTED TOGTHER
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.ROUTER_PKG.ALL;

ENTITY ROUTERS_5_AND_6 IS
	GENERIC(
		ROUTER5_ADDRESS : NETWORK_ADDR;
		ROUTER6_ADDRESS : NETWORK_ADDR
	);
	PORT(
		-- GLOBAL CLOCK AND RESET SIGNALS
        	CLK                 : IN STD_LOGIC;
        	RST                 : IN STD_LOGIC;
		-- HANDLING INPUT BUFFERS
		-- INPUT PORTS FOR ADJACENT ROUTERS
		-- ROUTER 5 
        	NORTH_DATA_IN_5     : IN FLIT;
        	SOUTH_DATA_IN_5     : IN FLIT;
        	WEST_DATA_IN_5      : IN FLIT;
		-- ROUTER 6 
        	NORTH_DATA_IN_6     : IN FLIT;
        	EAST_DATA_IN_6      : IN FLIT;
        	SOUTH_DATA_IN_6     : IN FLIT;
		-- PORTS FOR CHECKING CREDIT OUT OF ADJACENT BUFFERS
		-- ROUTER 5
        	NORTH_CREDIT_IN_5   : IN STD_LOGIC;
        	SOUTH_CREDIT_IN_5   : IN STD_LOGIC;
        	WEST_CREDIT_IN_5    : IN STD_LOGIC;
		-- ROUTER 6
        	NORTH_CREDIT_IN_6   : IN STD_LOGIC;
        	EAST_CREDIT_IN_6    : IN STD_LOGIC;
        	SOUTH_CREDIT_IN_6   : IN STD_LOGIC;
		-- WRITE REQUEST SIGNALS COMES FROM ADJACENT ROUTERS
		-- ROUTER 5
        	NORTH_WR_REQ_IN_5   : IN STD_LOGIC;
        	SOUTH_WR_REQ_IN_5   : IN STD_LOGIC;
        	WEST_WR_REQ_IN_5    : IN STD_LOGIC;
		-- ROUTER 6
        	NORTH_WR_REQ_IN_6   : IN STD_LOGIC;
        	EAST_WR_REQ_IN_6    : IN STD_LOGIC;
        	SOUTH_WR_REQ_IN_6   : IN STD_LOGIC;
		-- OUTPUT PORTS TO ADJACENT ROUTERS 
		-- ROUTER 5
		LOCAL_DATA_OUT_5    : OUT FLIT;
        	NORTH_DATA_OUT_5    : OUT FLIT;
        	SOUTH_DATA_OUT_5    : OUT FLIT;
        	WEST_DATA_OUT_5     : OUT FLIT;
		-- ROUTER 6
		LOCAL_DATA_OUT_6    : OUT FLIT;
        	NORTH_DATA_OUT_6    : OUT FLIT;
        	EAST_DATA_OUT_6     : OUT FLIT;
        	SOUTH_DATA_OUT_6    : OUT FLIT;
		-- ROUTER'S OUTPUT SIGNALS
		-- ROUTER 5
		LOCAL_CREDIT_OUT_5  : OUT STD_LOGIC;
        	NORTH_CREDIT_OUT_5  : OUT STD_LOGIC;
        	SOUTH_CREDIT_OUT_5  : OUT STD_LOGIC;
        	WEST_CREDIT_OUT_5   : OUT STD_LOGIC;
		-- ROUTER 6
		LOCAL_CREDIT_OUT_6  : OUT STD_LOGIC;
        	NORTH_CREDIT_OUT_6  : OUT STD_LOGIC;
        	EAST_CREDIT_OUT_6   : OUT STD_LOGIC;
        	SOUTH_CREDIT_OUT_6  : OUT STD_LOGIC;
		-- WRITE REQUEST SIGNALS TO ADJACENT ROUTERS
		-- ROUTER 5
        	NORTH_WR_REQ_OUT_5  : OUT STD_LOGIC;
        	SOUTH_WR_REQ_OUT_5  : OUT STD_LOGIC;
        	WEST_WR_REQ_OUT_5   : OUT STD_LOGIC;
		-- ROUTER 6
        	NORTH_WR_REQ_OUT_6  : OUT STD_LOGIC;
        	EAST_WR_REQ_OUT_6   : OUT STD_LOGIC;
        	SOUTH_WR_REQ_OUT_6  : OUT STD_LOGIC;
		-- IP CORE RELATED SIGNALS
		-- ROUTER 5
		FLIT_DEST_ADDR_TO_NI_5 : IN    NETWORK_ADDR;
		HEAD_OR_TAIL_5         : IN    STD_LOGIC;
        	VALID_TO_NI_5          : IN    STD_LOGIC;
		READY_FROM_NI_5        : OUT   STD_LOGIC;
		READY_TO_NI_5          : IN    STD_LOGIC;                                    
        	PAYLOAD_FORM_NI_5      : OUT   STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        	VALID_FROM_NI_5        : OUT   STD_LOGIC;
		-- ROUTER 6
		FLIT_DEST_ADDR_TO_NI_6 : IN    NETWORK_ADDR;
		HEAD_OR_TAIL_6         : IN    STD_LOGIC;
        	VALID_TO_NI_6          : IN    STD_LOGIC;
		READY_FROM_NI_6        : OUT   STD_LOGIC;
		READY_TO_NI_6          : IN    STD_LOGIC;                                    
        	PAYLOAD_FORM_NI_6      : OUT   STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        	VALID_FROM_NI_6        : OUT   STD_LOGIC
	);

END ENTITY ROUTERS_5_AND_6;

ARCHITECTURE STRUCT OF ROUTERS_5_AND_6 IS

-- COMPONENT DECLARATION
COMPONENT ROUTER 
	GENERIC(
		NODE_ADDRESS : NETWORK_ADDR
	);
	PORT(
		-- GLOBAL CLOCK AND RESET SIGNALS
        	CLK               : IN STD_LOGIC;
        	RST               : IN STD_LOGIC;
		-- HANDLING INPUT BUFFERS
		-- INPUT PORTS FOR ADJACENT ROUTERS
        	NORTH_DATA_IN     : IN FLIT;
        	EAST_DATA_IN      : IN FLIT;
        	SOUTH_DATA_IN     : IN FLIT;
        	WEST_DATA_IN      : IN FLIT;
		-- PORTS FOR CHECKING CREDIT OUT OF ADJACENT BUFFERS
        	NORTH_CREDIT_IN   : IN STD_LOGIC;
        	EAST_CREDIT_IN    : IN STD_LOGIC;
        	SOUTH_CREDIT_IN   : IN STD_LOGIC;
        	WEST_CREDIT_IN    : IN STD_LOGIC;
		-- WRITE REQUEST SIGNALS COMES FROM ADJACENT ROUTERS
        	NORTH_WR_REQ_IN   : IN STD_LOGIC;
        	EAST_WR_REQ_IN    : IN STD_LOGIC;
        	SOUTH_WR_REQ_IN   : IN STD_LOGIC;
        	WEST_WR_REQ_IN    : IN STD_LOGIC;
		-- OUTPUT PORTS TO ADJACENT ROUTERS 
		LOCAL_DATA_OUT    : OUT FLIT;
        	NORTH_DATA_OUT    : OUT FLIT;
        	EAST_DATA_OUT     : OUT FLIT;
        	SOUTH_DATA_OUT    : OUT FLIT;
        	WEST_DATA_OUT     : OUT FLIT;
		-- ROUTER'S OUTPUT SIGNALS
		LOCAL_CREDIT_OUT  : OUT STD_LOGIC;
        	NORTH_CREDIT_OUT  : OUT STD_LOGIC;
        	EAST_CREDIT_OUT   : OUT STD_LOGIC;
        	SOUTH_CREDIT_OUT  : OUT STD_LOGIC;
        	WEST_CREDIT_OUT   : OUT STD_LOGIC;
		-- WRITE REQUEST SIGNALS TO ADJACENT ROUTERS
        	NORTH_WR_REQ_OUT  : OUT STD_LOGIC;
        	EAST_WR_REQ_OUT   : OUT STD_LOGIC;
        	SOUTH_WR_REQ_OUT  : OUT STD_LOGIC;
        	WEST_WR_REQ_OUT   : OUT STD_LOGIC;
		-- IP CORE RELATED SIGNALS
		FLIT_DEST_ADDR_TO_NI : IN    NETWORK_ADDR;
		HEAD_OR_TAIL         : IN    STD_LOGIC;
        	VALID_TO_NI          : IN    STD_LOGIC;
		READY_FROM_NI        : OUT   STD_LOGIC;
		READY_TO_NI          : IN    STD_LOGIC;                                    
        	PAYLOAD_FORM_NI      : OUT   STD_LOGIC_VECTOR(ADDRESS_WIDTH - 1 DOWNTO 0);
        	VALID_FROM_NI        : OUT   STD_LOGIC
	);

END COMPONENT;

-- SIGNALS AND INTERCONNECTIONS

-- INPUT DATA OF BOTH ROUTERS
SIGNAL EAST_DATA_IN5, WEST_DATA_IN6 : FLIT;

-- OUTPUTS OF BOTH ROUTERS 
-- ROUTER 5
SIGNAL LDO5, NDO5, SDO5, WDO5 : FLIT;
-- ROUTER 6
SIGNAL LDO6, NDO6, EDO6, SDO6 : FLIT;

-- CREDIT IN OF BOTH ROUTERS
SIGNAL EAST_CREDIT_IN_5, WEST_CREDIT_IN_6 : STD_LOGIC;

-- CREDIT OUT OF BOTH ROUTERS
-- ROUTER 5
SIGNAL LCO5, NCO5, SCO5, WCO5 : STD_LOGIC;
-- ROUTER 6
SIGNAL LCO6, NCO6, ECO6, SCO6 : STD_LOGIC;

-- WRITE REQUEST IN OF BOTH ROUTERS
SIGNAL EAST_WR_REQ_IN_5, WEST_WR_REQ_IN_6 : STD_LOGIC;

-- WRITE REQUEST OUT OF BOTH ROUTERS
-- ROUTER 5
SIGNAL NWRO5, SWRO5, WWRO5 : STD_LOGIC;
-- ROUTER 6
SIGNAL NWRO6, EWRO6, SWRO6 : STD_LOGIC;

-- IP CORE RELATED SIGNALS
SIGNAL RFNI5, RFNI6, VFNI5, VFNI6 : STD_LOGIC;
SIGNAL PFNI5, PFNI6 : NETWORK_ADDR;

BEGIN

-- COMPONENT INSTATIATION
-- ROUTER 5
ROUTER5 : ROUTER 
	GENERIC MAP(
		NODE_ADDRESS      => ROUTER5_ADDRESS
	)
	PORT MAP(
		-- GLOBAL CLOCK AND RESET SIGNALS
        	CLK               => CLK,
        	RST               => RST,
		-- HANDLING INPUT BUFFERS
		-- INPUT PORTS FOR ADJACENT ROUTERS
        	NORTH_DATA_IN     => NORTH_DATA_IN_5,
        	EAST_DATA_IN      => EAST_DATA_IN5,
        	SOUTH_DATA_IN     => SOUTH_DATA_IN_5,
        	WEST_DATA_IN      => WEST_DATA_IN_5,
		-- PORTS FOR CHECKING CREDIT OUT OF ADJACENT BUFFERS
        	NORTH_CREDIT_IN   => NORTH_CREDIT_IN_5,
        	EAST_CREDIT_IN    => EAST_CREDIT_IN_5,
        	SOUTH_CREDIT_IN   => SOUTH_CREDIT_IN_5,
        	WEST_CREDIT_IN    => WEST_CREDIT_IN_5,
		-- WRITE REQUEST SIGNALS COMES FROM ADJACENT ROUTERS
        	NORTH_WR_REQ_IN   => NORTH_WR_REQ_IN_5,
        	EAST_WR_REQ_IN    => EAST_WR_REQ_IN_5,
        	SOUTH_WR_REQ_IN   => SOUTH_WR_REQ_IN_5,
        	WEST_WR_REQ_IN    => WEST_WR_REQ_IN_5,
		-- OUTPUT PORTS TO ADJACENT ROUTERS 
		LOCAL_DATA_OUT    => LDO5,
        	NORTH_DATA_OUT    => NDO5,
        	EAST_DATA_OUT     => WEST_DATA_IN6,
        	SOUTH_DATA_OUT    => SDO5,
        	WEST_DATA_OUT     => WDO5,
		-- ROUTER'S OUTPUT SIGNALS
		LOCAL_CREDIT_OUT  => LCO5,
        	NORTH_CREDIT_OUT  => NCO5,
        	EAST_CREDIT_OUT   => WEST_CREDIT_IN_6,
        	SOUTH_CREDIT_OUT  => SCO5,
        	WEST_CREDIT_OUT   => WCO5,
		-- WRITE REQUEST SIGNALS TO ADJACENT ROUTERS
        	NORTH_WR_REQ_OUT  => NWRO5,
        	EAST_WR_REQ_OUT   => WEST_WR_REQ_IN_6,
        	SOUTH_WR_REQ_OUT  => SWRO5,
        	WEST_WR_REQ_OUT   => WWRO5,
		-- IP CORE RELATED SIGNALS
		FLIT_DEST_ADDR_TO_NI => FLIT_DEST_ADDR_TO_NI_5,
		HEAD_OR_TAIL         => HEAD_OR_TAIL_5,
        	VALID_TO_NI          => VALID_TO_NI_5,
		READY_FROM_NI        => RFNI5,
		READY_TO_NI          => READY_TO_NI_5,                                    
        	PAYLOAD_FORM_NI      => PFNI5,
        	VALID_FROM_NI        => VFNI5
	);

-- ROUTER 6
ROUTER6 : ROUTER 
	GENERIC MAP(
		NODE_ADDRESS      => ROUTER6_ADDRESS
	)
	PORT MAP(
		-- GLOBAL CLOCK AND RESET SIGNALS
        	CLK               => CLK,
        	RST               => RST,
		-- HANDLING INPUT BUFFERS
		-- INPUT PORTS FOR ADJACENT ROUTERS
        	NORTH_DATA_IN     => NORTH_DATA_IN_6,
        	EAST_DATA_IN      => EAST_DATA_IN_6,
        	SOUTH_DATA_IN     => SOUTH_DATA_IN_6,
        	WEST_DATA_IN      => WEST_DATA_IN6,
		-- PORTS FOR CHECKING CREDIT OUT OF ADJACENT BUFFERS
        	NORTH_CREDIT_IN   => NORTH_CREDIT_IN_6,
        	EAST_CREDIT_IN    => EAST_CREDIT_IN_6,
        	SOUTH_CREDIT_IN   => SOUTH_CREDIT_IN_6,
        	WEST_CREDIT_IN    => WEST_CREDIT_IN_6,
		-- WRITE REQUEST SIGNALS COMES FROM ADJACENT ROUTERS
        	NORTH_WR_REQ_IN   => NORTH_WR_REQ_IN_6,
        	EAST_WR_REQ_IN    => EAST_WR_REQ_IN_6,
        	SOUTH_WR_REQ_IN   => SOUTH_WR_REQ_IN_6,
        	WEST_WR_REQ_IN    => WEST_WR_REQ_IN_6,
		-- OUTPUT PORTS TO ADJACENT ROUTERS 
		LOCAL_DATA_OUT    => LDO6,
        	NORTH_DATA_OUT    => NDO6,
        	EAST_DATA_OUT     => EDO6,
        	SOUTH_DATA_OUT    => SDO6,
        	WEST_DATA_OUT     => EAST_DATA_IN5,
		-- ROUTER'S OUTPUT SIGNALS
		LOCAL_CREDIT_OUT  => LCO6,
        	NORTH_CREDIT_OUT  => NCO6,
        	EAST_CREDIT_OUT   => ECO6,
        	SOUTH_CREDIT_OUT  => SCO6,
        	WEST_CREDIT_OUT   => EAST_CREDIT_IN_5,
		-- WRITE REQUEST SIGNALS TO ADJACENT ROUTERS
        	NORTH_WR_REQ_OUT  => NWRO6,
        	EAST_WR_REQ_OUT   => EWRO6,
        	SOUTH_WR_REQ_OUT  => SWRO6,
        	WEST_WR_REQ_OUT   => EAST_WR_REQ_IN_5,
		-- IP CORE RELATED SIGNALS
		FLIT_DEST_ADDR_TO_NI => FLIT_DEST_ADDR_TO_NI_6,
		HEAD_OR_TAIL         => HEAD_OR_TAIL_6,
        	VALID_TO_NI          => VALID_TO_NI_6,
		READY_FROM_NI        => RFNI6,
		READY_TO_NI          => READY_TO_NI_6,                                    
        	PAYLOAD_FORM_NI      => PFNI6,
        	VALID_FROM_NI        => VFNI6
	);

	-- CREDIT OUTS
	-- ROUTER 5
	LOCAL_CREDIT_OUT_5  <= LCO5;
        NORTH_CREDIT_OUT_5  <= NCO5;
        SOUTH_CREDIT_OUT_5  <= SCO5;
        WEST_CREDIT_OUT_5   <= WCO5;
	-- ROUTER 6
	LOCAL_CREDIT_OUT_6  <= LCO6;
        NORTH_CREDIT_OUT_6  <= NCO6;
        EAST_CREDIT_OUT_6   <= ECO6;
        SOUTH_CREDIT_OUT_6  <= SCO6;
	-- WRITE REQUEST OUT
	-- ROUTER 5
        NORTH_WR_REQ_OUT_5  <= NWRO5;
        SOUTH_WR_REQ_OUT_5  <= SWRO5;
        WEST_WR_REQ_OUT_5   <= WWRO5;
	-- ROUTER 6
        NORTH_WR_REQ_OUT_6  <= NWRO6;
        EAST_WR_REQ_OUT_6   <= EWRO6;
        SOUTH_WR_REQ_OUT_6  <= SWRO6;
	-- OUTPUTS ADJACENT ROUTERS 
	-- ROUTER 5
	LOCAL_DATA_OUT_5    <= LDO5;
        NORTH_DATA_OUT_5    <= NDO5;
        SOUTH_DATA_OUT_5    <= SDO5;
        WEST_DATA_OUT_5     <= WDO5;
	-- ROUTER 6
	LOCAL_DATA_OUT_6    <= LDO6;
        NORTH_DATA_OUT_6    <= NDO6;
        EAST_DATA_OUT_6     <= EDO6;
        SOUTH_DATA_OUT_6    <= SDO6;

	-- IP CORE 
	--ROUTER 5
	READY_FROM_NI_5     <= RFNI5;
	PAYLOAD_FORM_NI_5   <= PFNI5;
	VALID_FROM_NI_5     <= VFNI5;
	--ROUTER 6
	READY_FROM_NI_6     <= RFNI6;
	PAYLOAD_FORM_NI_6   <= PFNI6;
	VALID_FROM_NI_6     <= VFNI6;

END ARCHITECTURE;
